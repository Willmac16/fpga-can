// Can2040 will hit 1Mbit/s == 1 microsecond nominal bit time
// Alchitry Clock is 100 MHz == 0.01 microseconds per clock
// 100 quanta per bit time

`timescale 10 ns / 1 ps

module recieve_tb;
    reg updated_sample, rx, stuff_error;

    wire [63:0] msg;
    wire [28:0] msg_id;
    wire rtr, extended, bus_idle, FORM_ERROR, OVERLOAD_ERROR, fire_an_ack, msg_fresh;

    reg next_bit, clear_crc, update_crc;

    wire [14:0] crc;

    message_reciever reciever (.updated_sample(updated_sample), .stuff_error(stuff_error), .rx(rx), .msg_id(msg_id), .rtr(rtr), .extended(extended), .msg(msg), .bus_idle(bus_idle), .stuff_bypass(stuff_bypass), .FORM_ERROR(FORM_ERROR), .OVERLOAD_ERROR(OVERLOAD_ERROR), .fire_an_ack(fire_an_ack), .msg_fresh(msg_fresh));
    crc_step_machine crcsm (.next_bit(next_bit), .clear_crc(clear_crc), .update_crc(update_crc), .crc(crc));

    reg [163:0] test_stream;
    integer i;

    initial begin
        $dumpfile("can.lx2");
        $dumpvars(0, reciever);
        $dumpvars(0, test_stream);
        $dumpvars(0, crcsm);

        // Init
        stuff_error <= 0;
        updated_sample <= 0;

        // Valid MSG
        test_stream[63] <= 1; // SOF
        test_stream[62:52] <= 11'b01100110011; // ID
        test_stream[51] <= 1; // RTR
        test_stream[50:49] <= 2'b11; // Reserved
        test_stream[48:45] <= 4'd0; // DLC

        test_stream[44:30] <= 15'd0; // CRC
        test_stream[29] <= 1'b0; // CRC Delim

        test_stream[28] <= 1'b1; // ACK
        test_stream[27] <= 1'b0; // ACK Delim

        test_stream[26:20] <= 7'b0000000; // EOF
        test_stream[19:0] <= 0;

        clear_crc <= 1;
        #1;

        clear_crc <= 0;
        #1;

        for (i = 63; i >= 45; i = i - 1) begin
            next_bit <= test_stream[i];
            update_crc <= 1;
            #0.01;
            update_crc <= 0;
            #0.01;
        end

        test_stream[44:30] <= crc;

        #1;

        for (i = 63; i >= 0; i = i - 1) begin
            rx = test_stream[i];
            updated_sample = 1;
            #1;
            updated_sample = 0;
            #1;
        end

        // Valid Form, but invalid CRC
        test_stream[44:30] <= crc ^ 15'b011000101010011;
        #1;

        for (i = 63; i >= 0; i = i - 1) begin
            rx = test_stream[i];
            updated_sample = 1;
            #1;
            updated_sample = 0;
            #1;
        end

        // Msg with data
        test_stream[163] <= 1; // SOF
        test_stream[162:152] <= 11'b10001010101; // ID
        test_stream[151] <= 1; // RTR
        test_stream[150:149] <= 2'b11; // Reserved
        test_stream[148:145] <= 4'b1000; // DLC
        test_stream[144:81] <= 64'hd3359da81bd963e5; // Data

        test_stream[80:66] <= 15'd0; // CRC
        test_stream[65] <= 1'b0; // CRC Delim

        test_stream[64] <= 1'b1; // ACK
        test_stream[63] <= 1'b0; // ACK Delim

        test_stream[62:55] <= 7'b0000000; // EOF
        test_stream[54:0] <= 0;

        clear_crc <= 1;
        #1;

        clear_crc <= 0;
        #1;

        for (i = 163; i >= 81; i = i - 1) begin
            next_bit <= test_stream[i];
            update_crc <= 1;
            #0.01;
            update_crc <= 0;
            #0.01;
        end

        test_stream[80:66] <= crc;

        #1;

        for (i = 163; i >= 0; i = i - 1) begin
            rx = test_stream[i];
            updated_sample = 1;
            #1;
            updated_sample = 0;
            #1;
        end

        // Msg with data
        // Invalid CRC
        test_stream[163] <= 1; // SOF
        test_stream[162:152] <= 11'b10001010101; // ID
        test_stream[151] <= 1; // RTR
        test_stream[150:149] <= 2'b11; // Reserved
        test_stream[148:145] <= 4'b1000; // DLC
        test_stream[144:81] <= 64'hd3359da81bd963e5; // Data

        test_stream[80:66] <= 15'd0; // CRC
        test_stream[65] <= 1'b0; // CRC Delim

        test_stream[64] <= 1'b1; // ACK
        test_stream[63] <= 1'b0; // ACK Delim

        test_stream[62:55] <= 7'b0000000; // EOF
        test_stream[54:0] <= 0;

        clear_crc <= 1;
        #1;

        clear_crc <= 0;
        #1;

        for (i = 163; i >= 81; i = i - 1) begin
            next_bit <= test_stream[i];
            update_crc <= 1;
            #0.01;
            update_crc <= 0;
            #0.01;
        end

        test_stream[80:66] <= ~crc;

        #1;

        for (i = 163; i >= 0; i = i - 1) begin
            rx = test_stream[i];
            updated_sample = 1;
            #1;
            updated_sample = 0;
            #1;
        end

        // Extended ID Msg with data
        test_stream[163] <= 1; // SOF
        test_stream[162:152] <= ~11'b10001010101; // Base ID
        test_stream[151] <= 0; // SRR
        test_stream[150] <= 0; // IDE
        test_stream[149:132] <= 18'b100010101010101010; // Extended ID
        test_stream[131] <= 1; // RTR
        test_stream[130:129] <= 2'b11; // Reserved
        test_stream[128:125] <= 4'b1000; // DLC
        test_stream[124:61] <= 64'hd3359da81bd963e5 ^ 64'b1010101010101010101010101010101010101010101010101010101010101010; // Datas
        test_stream[45] <= 1'b0; // CRC Delim

        test_stream[44] <= 1'b1; // ACK
        test_stream[43] <= 1'b0; // ACK Delim

        test_stream[42:35] <= 7'b0000000; // EOF
        test_stream[34:0] <= 0;

        clear_crc <= 1;
        #1;

        clear_crc <= 0;
        #1;

        for (i = 163; i >= 61; i = i - 1) begin
            next_bit <= test_stream[i];
            update_crc <= 1;
            #0.01;
            update_crc <= 0;
            #0.01;
        end

        test_stream[60:46] <= crc;

        #1;

        for (i = 163; i >= 0; i = i - 1) begin
            rx = test_stream[i];
            updated_sample = 1;
            #1;
            updated_sample = 0;
            #1;
        end

        // High CRC Delim
        test_stream[45] <= 1'b1; // CRC Delim

        #1;

        for (i = 163; i >= 0; i = i - 1) begin
            rx = test_stream[i];
            updated_sample = 1;
            #1;
            updated_sample = 0;
            #1;
        end

        // High Ack Delim
        test_stream[43] <= 1'b1; // CRC Delim

        #1;

        for (i = 163; i >= 0; i = i - 1) begin
            rx = test_stream[i];
            updated_sample = 1;
            #1;
            updated_sample = 0;
            #1;
        end


    end
endmodule

module crc_tb;
    reg next_bit, clear_crc, update_crc;
    wire [14:0] crc;
    reg [63:0] test_stream;

    integer i;

    crc_step_machine crcsm (.next_bit(next_bit), .clear_crc(clear_crc), .update_crc(update_crc), .crc(crc));
    initial begin
        $dumpfile("can.lx2");
        $dumpvars(0, test_stream);
        $dumpvars(0, crcsm);

        // Init
        clear_crc <= 1;
        #1;
        clear_crc <= 0;
        #1;

        // Test Stream
        test_stream = 64'hd3359da81bd963e5;
        for (i = 63; i >= 0; i = i - 1) begin
            next_bit <= test_stream[i];
            update_crc <= 1;
            #1;
            update_crc <= 0;
            #1;
        end

        $display("Data: %h", test_stream);
        $display("CRC: %h", crc);
    end
endmodule

module txp_tb;
    reg next_bit, updated_sample, rx_updated_sample, stuff_bypass, rx;
    wire tx, bit_advance, stuff_error, out_bit, doorbell;
    reg sync_tick;

    reg [23:0] txp_test_stream;
    reg [23:0] txp_out_stream;

    integer i;

    tx_pipeline txp (.tx(tx), .updated_sample(updated_sample), .next_bit(next_bit), .bit_advance(bit_advance), .stuff_bypass(stuff_bypass));
    rx_pipeline rxp (.rx(rx), .updated_sample(rx_updated_sample), .updated_bit(doorbell), .next_bit(out_bit), .stuff_error(stuff_error), .stuff_bypass(stuff_bypass));

    initial begin
        $dumpfile("can.lx2");
        $dumpvars(0, txp_test_stream);
        $dumpvars(0, txp_out_stream);
        $dumpvars(0, txp);
        $dumpvars(0, rxp);

        // Init
        stuff_bypass <= 1;
        #1
        stuff_bypass <= 0;
        updated_sample <= 0;
        rx_updated_sample <= 0;
        #1;

        // Stream without the need for stuff
        txp_test_stream = 24'b100100100100100100100100;
        i = 23;
        while (i >= 0) begin
            next_bit <= txp_test_stream[i];
            updated_sample <= 1;
            #1;
            rx <= tx;
            rx_updated_sample <= 1;
            if (bit_advance) begin
                i = i - 1;
            end

            #1
            if (doorbell) begin
                txp_out_stream <= {txp_out_stream[22:0], out_bit};
            end
            #1;
            updated_sample <= 0;
            rx_updated_sample <= 0;
            #1;
        end

        stuff_bypass <= 1;
        #1;
        stuff_bypass <= 0;

        // Stream with stuffing
        txp_test_stream = 24'b100000000011111111100000;
        i = 23;
        #1;
        while (i >= 0) begin
            next_bit <= txp_test_stream[i];
            updated_sample <= 1;
            #1;
            rx <= tx;
            rx_updated_sample <= 1;
            if (bit_advance) begin
                i = i - 1;
            end

            #1
            if (doorbell) begin
                txp_out_stream <= {txp_out_stream[22:0], out_bit};
            end
            #1;
            updated_sample <= 0;
            rx_updated_sample <= 0;
            #1;
        end
    end
endmodule

module rxp_tb;
    reg rx, updated_sample, stuff_bypass;
    wire updated_bit, next_bit, stuff_error;

    reg [23:0] test_stream;
    reg [23:0] out_stream;

    integer i;

    rx_pipeline rxp (.rx(rx), .updated_sample(updated_sample), .updated_bit(updated_bit), .next_bit(next_bit), .stuff_error(stuff_error), .stuff_bypass(stuff_bypass));

    initial begin
        $dumpfile("can.lx2");
        $dumpvars(0, test_stream);
        $dumpvars(0, out_stream);
        $dumpvars(0, rxp);

        // Init
        stuff_bypass <= 1;
        #1
        stuff_bypass <= 0;
        rx <= 0;
        updated_sample <= 0;
        #1;

        // Valid Data Stream without Stuff
        test_stream = 24'b100100100100100100100100;
        for (i = 23; i >= 0; i = i - 1) begin
            rx <= test_stream[i];
            #1;
            updated_sample <= 1;
            #1;
            if (updated_bit) begin
                out_stream <= {next_bit, out_stream[23:1]};
            end
            updated_sample <= 0;
        end

        stuff_bypass <= 1;
        #1;
        stuff_bypass <= 0;

        // Valid Data Stream with Stuff
        test_stream = 24'b100000100011111011110010;
        #1
        for (i = 23; i >= 0; i = i - 1) begin
            rx <= test_stream[i];
            #1;
            updated_sample <= 1;
            #1;
            if (updated_bit) begin
                out_stream <= {next_bit, out_stream[23:1]};
            end
            updated_sample <= 0;
        end

        stuff_bypass <= 1;
        #1;
        for (i = 23; i >= 0; i = i - 1) begin
            rx <= test_stream[i];
            #1;
            updated_sample <= 1;
            #1;
            if (updated_bit) begin
                out_stream <= {next_bit, out_stream[23:1]};
            end
            updated_sample <= 0;
        end

        stuff_bypass <= 0;
        #1;

        // Stuff Error Test
        test_stream = 24'b100000000011111111100000;
        #1
        for (i = 23; i >= 0; i = i - 1) begin
            rx <= test_stream[i];
            #1;
            updated_sample <= 1;
            #1;
            if (updated_bit) begin
                out_stream <= {next_bit, out_stream[23:1]};
            end
            updated_sample <= 0;
        end
    end
endmodule

module ssm_tb;
    reg rx_raw, clk, bus_idle;
    wire rx;
    reg [6:0] RJW;

    reg [123:0] can_test;

    always @(rx) begin
        bus_idle = 0;
    end

    sync_sample_machine ssm (.rx_raw(rx_raw), .clk(clk), .RJW(RJW), .bus_idle(bus_idle), .rx(rx));
    initial begin
        can_test[123] = 1;
        can_test[122:112] = 11'b1001001001;
        can_test[111:110] = 2'b00; // SRR & IDE
        can_test[109:92] = 18'b100100100100100100; // Extended ID
        can_test[91:89] = 3'b111; // RTR & R0 & R1
        can_test[88:85] = 4'b0001; // DLC
        can_test[84:77] = 8'b01010101; // Data Byte
        can_test[76:62] = 15'b100100100100100; // CRC
        can_test[61:52] = 10'b0100000000; // Delims, ACK & EOF
        can_test[51:0] = 52'b0; // Bus Idle



        // $dumpfile("can.vcd");
        $dumpvars(0, ssm);
        clk = 0;
        RJW = 1;
        bus_idle = 1;
        rx_raw = 0;
        #1;

        for (integer i = 123; i > 0; i = i - 1) begin
            rx_raw = can_test[i];
            for (integer i = 0; i < 100; i = i + 1) begin
                clk = 1;
                #0.45;
                clk = 0;
                #0.45;
            end
        end


    end
endmodule
